library IEEE;
use IEEE.STD_LOGIC_1164.all;

package ReactTimePack is
 
  constant DISABLE_PAT : std_logic_vector(6 downto 0) := "1111111";
  constant HYPHEN_PAT  : std_logic_vector(6 downto 0) := "0111111";
  constant DISP_C      : std_logic_vector(6 downto 0) := "1000110";
  constant DISP_O      : std_logic_vector(6 downto 0) := "1000000";
  constant DISP_N      : std_logic_vector(6 downto 0) := "0101011";
  constant DISP_F      : std_logic_vector(6 downto 0) := "0001110";
  constant DISP_T      : std_logic_vector(6 downto 0) := "0000111";
  constant DISP_E      : std_logic_vector(6 downto 0) := "0000110";
  constant DISP_S      : std_logic_vector(6 downto 0) := "0010010";
  
end package ReactTimePack;
 

package body ReactTimePack is
end package body ReactTimePack;

